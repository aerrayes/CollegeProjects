module muxx ( s , w , f);
input [2:0] s ;
input [7:0] w ;
output F;

