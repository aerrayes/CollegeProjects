module Decrement (a,cin,f,cout);
	input a,cin;
	output f,cout;
	Full_adder x (a,1,cin,f,cout);
endmodule
